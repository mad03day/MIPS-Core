`timescale 1 ns / 10 ps

module testbench;

reg i_clk_r, i_rst_n_r;
parameter period = 100;

mips testbench(.clk(i_clk_r), .reset(i_rst_n_r));

initial
begin
#8000 $finish;
end 
initial
begin
i_clk_r = 0;
forever#(period/2) i_clk_r = ~i_clk_r;
end
initial
begin
i_rst_n_r = 0;
#125 i_rst_n_r = 1;
end
endmodule
 //                              100 01000 00011 00000 100000
//   hex 00881820 bin 000000 00100 01000 00011 00000 100000 000000/op 00100/rs-r4 01000/rt-r8 00011/rd-3 100000 /ifunc Add (00000000100010000001100000100000)
//                               100 01000 00011 00000 100100
//   hex 00881824 bin 000000 00100 01000 00011 00000 100100 000000/op 00100/rs-r4 01000/rt-r8 00011/rd-3 100100 /ifunc AND (00000000100010000001100000100100)
//   hex 2025003F bin 001000 00001 11100 0000000000111111     001000/op(addi)   00001/rs-r1  11100/rd-r28  00000 00000 111111 imm
//   hex 8CE20000 bin 100011 00111 00010 0000000000000000     100011/op(lw)   00111/rs-r7    00010/rd-r2 0000000000000000 imm

//                      101011 00111 00100 0000 0000 0000 0000
//   hex ACE40000 bin 101011 00111 00100 0000000000000000     101011/op(sw)   00111/rs-r7    00100/rd-r4 0000000000000000 imm (10101100111000000000000000000000)
//   hex 10000001 bin 000100 00000 00000 00000 00000 000001     000100/op(beq)   0000000000   00000 00000 000001 ofset
//   hex 08000000 bin 000010 00000 00000 00000 00000 000100     000010/op(j)   00000 00000 00000 00000 000000 imm